// megafunction wizard: %LPM_DIVIDE%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: LPM_DIVIDE 

// ============================================================
// File Name: divide_9d7.v
// Megafunction Name(s):
// 			LPM_DIVIDE
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 10.1 Build 197 01/19/2011 SP 1 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module divide_9d7 (
	denom,
	numer,
	quotient,
	remain);

	input	[6:0]  denom;
	input	[8:0]  numer;
	output	[8:0]  quotient;
	output	[6:0]  remain;

	wire [8:0] sub_wire0;
	wire [6:0] sub_wire1;
	wire [8:0] quotient = sub_wire0[8:0];
	wire [6:0] remain = sub_wire1[6:0];

	lpm_divide	LPM_DIVIDE_component (
				.denom (denom),
				.numer (numer),
				.quotient (sub_wire0),
				.remain (sub_wire1),
				.aclr (1'b0),
				.clken (1'b1),
				.clock (1'b0));
	defparam
		LPM_DIVIDE_component.lpm_drepresentation = "UNSIGNED",
		LPM_DIVIDE_component.lpm_hint = "MAXIMIZE_SPEED=6,LPM_REMAINDERPOSITIVE=TRUE",
		LPM_DIVIDE_component.lpm_nrepresentation = "UNSIGNED",
		LPM_DIVIDE_component.lpm_type = "LPM_DIVIDE",
		LPM_DIVIDE_component.lpm_widthd = 7,
		LPM_DIVIDE_component.lpm_widthn = 9;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: PRIVATE: PRIVATE_LPM_REMAINDERPOSITIVE STRING "TRUE"
// Retrieval info: PRIVATE: PRIVATE_MAXIMIZE_SPEED NUMERIC "6"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: USING_PIPELINE NUMERIC "0"
// Retrieval info: PRIVATE: VERSION_NUMBER NUMERIC "2"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_DREPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: LPM_HINT STRING "MAXIMIZE_SPEED=6,LPM_REMAINDERPOSITIVE=TRUE"
// Retrieval info: CONSTANT: LPM_NREPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_DIVIDE"
// Retrieval info: CONSTANT: LPM_WIDTHD NUMERIC "7"
// Retrieval info: CONSTANT: LPM_WIDTHN NUMERIC "9"
// Retrieval info: USED_PORT: denom 0 0 7 0 INPUT NODEFVAL "denom[6..0]"
// Retrieval info: USED_PORT: numer 0 0 9 0 INPUT NODEFVAL "numer[8..0]"
// Retrieval info: USED_PORT: quotient 0 0 9 0 OUTPUT NODEFVAL "quotient[8..0]"
// Retrieval info: USED_PORT: remain 0 0 7 0 OUTPUT NODEFVAL "remain[6..0]"
// Retrieval info: CONNECT: @denom 0 0 7 0 denom 0 0 7 0
// Retrieval info: CONNECT: @numer 0 0 9 0 numer 0 0 9 0
// Retrieval info: CONNECT: quotient 0 0 9 0 @quotient 0 0 9 0
// Retrieval info: CONNECT: remain 0 0 7 0 @remain 0 0 7 0
// Retrieval info: GEN_FILE: TYPE_NORMAL divide_9d7.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL divide_9d7.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL divide_9d7.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL divide_9d7.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL divide_9d7_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL divide_9d7_bb.v FALSE
// Retrieval info: LIB_FILE: lpm
